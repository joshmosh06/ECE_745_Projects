//------------------------------------------------------------------------------
//
//  Description: I2c Package file that includes all files for the i2c package
//
//
//  Joshua Hofmann
//  North Carolina State University
//  3/9/2020
//  Built with ModelSim 10.6c
//------------------------------------------------------------------------------
package i2c_pkg;
	import ncsu_pkg::*;
	`include "src/i2c_typedefs.svh"
	`include "src/i2c_transaction.svh"
	`include "src/i2c_configuration.svh"
	`include "src/i2c_driver.svh"
	`include "src/i2c_monitor.svh"
	`include "src/i2c_agent.svh"


endpackage
