//I2cmb_env_pkg.sv file