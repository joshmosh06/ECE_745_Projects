//------------------------------------------------------------------------------
//
//  Description: wb configuration class
//
//
//  Joshua Hofmann
//  North Carolina State University
//  3/9/2020
//  Built with ModelSim 10.6c
//------------------------------------------------------------------------------
class wb_configuration extends ncsu_configuration;
  rand bit [5:0] min_delay;				//Randomized min/max Response Delay from slave
  rand bit [5:0] max_delay;
  rand bit       sop_eop_polarity;		//Randomized idk
  bit            enable;				//Enable slave
  bit            collect_coverage;		//Enable Coverage functionality
  //Min delay must be less than Max delay
constraint delay_range_c { min_delay < max_delay; }

covergroup wb_configuration_cg;
  	option.per_instance = 1;
    option.name = name;
  	coverpoint min_delay;
  	coverpoint max_delay;
  	coverpoint sop_eop_polarity;
  endgroup

  function void sample_coverage();
  	wb_configuration_cg.sample();
  endfunction
  
  function new(string name=""); 
    super.new(name);
    wb_configuration_cg = new;
  endfunction

  virtual function string convert2string();
     return {super.convert2string};
  endfunction

endclass : wb_configuration